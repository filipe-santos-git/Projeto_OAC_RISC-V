`timescale 1ns / 1ps

module Controller (
    //Input
    input logic [6:0] Opcode,
    //7-bit opcode field from the instruction

    //Outputs
    output logic ALUSrc,
    //0: The second ALU operand comes from the second register file output (Read data 2); 
    //1: The second ALU operand is the sign-extended, lower 16 bits of the instruction.
    output logic MemtoReg,
    //0: The value fed to the register Write data input comes from the ALU.
    //1: The value fed to the register Write data input comes from the data memory.
    output logic RegWrite, //The register on the Write register input is written with the value on the Write data input 
    output logic MemRead,  //Data memory contents designated by the address input are put on the Read data output
    output logic MemWrite, //Data memory contents designated by the address input are replaced by the value on the Write data input.
    output logic JalrSel, //1: BrPC = RD_One + ($signed(Imm)); 0: BrPC = (Branch_Sel) ? PC_Imm : 32'b0
    output logic jal_signal, //1: WB_Data = D.Pc_Four; 0: (D.lui_signal) ? D.ImmG : WrmuxSrc
    output logic lui_signal, //1: D.ImmG; 0: WrmuxSrc
    output logic [1:0] ALUOp,  //00: LW/SW; 01:Branch; 10: Rtype
    output logic Branch  //0: branch is not taken; 1: branch is taken
);

  logic [6:0] I_TYPE, R_TYPE, U_TYPE, LW, SW, BR, JAL, JALR, HALT;

  assign I_TYPE = 7'b0010011;   //addi,slti,slli,srli,srai
  assign R_TYPE = 7'b0110011;   //add,and,slt
  assign U_TYPE = 7'b0110111;   //lui
  assign LW     = 7'b0000011;   //lw
  assign SW     = 7'b0100011;   //sw
  assign BR     = 7'b1100011;   //beq,bne,blt,bge
  assign JAL    = 7'b1101111;   //jal
  assign JALR   = 7'b1100111;   //jalr
  assign HALT   = 7'b1111111;   //halt

  assign ALUSrc = (Opcode == LW || Opcode == SW || Opcode == I_TYPE || Opcode == JAL || Opcode == JALR);
  assign MemtoReg = (Opcode == LW);
  assign RegWrite = (Opcode == R_TYPE || Opcode == LW || Opcode == I_TYPE || Opcode == JAL || Opcode == JALR || Opcode == U_TYPE);
  assign MemRead = (Opcode == LW);
  assign MemWrite = (Opcode == SW);
  assign ALUOp[0] = (Opcode == BR || Opcode == JAL || Opcode == JALR);
  assign ALUOp[1] = (Opcode == R_TYPE || Opcode == I_TYPE || Opcode == JAL || Opcode == JALR);
  assign Branch = (Opcode == BR || Opcode == JAL || Opcode == JALR);
  assign JalrSel = (Opcode == JALR);
  assign jal_signal = (Opcode == JAL || Opcode == JALR);
  assign lui_signal = (Opcode == U_TYPE);
endmodule
